* Spice description of inversor_novo
* Spice driver version 270587057
* Date ( dd/mm/yyyy hh:mm:ss ): 26/05/2014 at 15:43:10

* INTERF a vdd vss y 


.subckt inversor_novo 1 2 4 3 
* NET 1 = a
* NET 2 = vdd
* NET 3 = y
* NET 4 = vss
Mtr_00002 2 1 3 2 tp L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00001 4 1 3 4 tn L=1U W=1U AS=2P AD=2P PS=6U PD=6U 
C4 1 4 1.697e-14
C3 2 4 9.03e-15
C2 3 4 1.003e-14
C1 4 4 9.03e-15
.ends inversor_novo


* Spice description of somador_1bit_genlib_ocp_1_rows_roteado
* Spice driver version 270587057
* Date ( dd/mm/yyyy hh:mm:ss ): 18/11/2014 at 15:29:32

* INTERF a b c r s vdd vss 


.subckt somador_1bit_genlib_ocp_1_rows_roteado 62 46 53 58 39 64 23 
* NET 23 = vss
* NET 24 = sinv10
* NET 25 = snand12
* NET 26 = snand10
* NET 27 = snand9
* NET 28 = snand8
* NET 29 = snand7
* NET 30 = sinv6
* NET 31 = sinv5
* NET 32 = snand6
* NET 33 = sinv7
* NET 34 = sinv9
* NET 35 = sinv8
* NET 36 = sinv1
* NET 37 = sinv4
* NET 38 = snand5
* NET 39 = s
* NET 40 = snand4
* NET 41 = snand21
* NET 42 = snand3
* NET 43 = snand16
* NET 44 = snand20
* NET 45 = sinv3
* NET 46 = b
* NET 47 = snand2
* NET 48 = snand15
* NET 49 = sinv13
* NET 50 = snand19
* NET 51 = snand14
* NET 52 = sinv12
* NET 53 = c
* NET 54 = snand18
* NET 55 = sinv2
* NET 56 = sinv15
* NET 57 = snand1
* NET 58 = r
* NET 59 = snand13
* NET 60 = sinv14
* NET 61 = sinv11
* NET 62 = a
* NET 63 = snand17
* NET 64 = vdd
Mtr_00118 63 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 64 61 63 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 61 59 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 58 60 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 64 56 58 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 57 55 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 64 53 57 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 54 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 64 52 54 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 52 51 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 50 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 64 49 50 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 49 48 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 47 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 64 45 47 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 60 44 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 44 43 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 64 63 44 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 42 55 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 64 45 42 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 56 41 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 40 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 64 53 40 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 41 54 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 64 50 41 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 38 36 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 64 37 38 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 39 35 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 64 34 39 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 33 40 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 32 36 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 64 31 32 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 36 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 29 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 64 30 29 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 30 42 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 28 62 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 64 33 28 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 31 47 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 27 38 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 64 32 27 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 26 29 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 64 28 26 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 37 57 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 45 53 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 25 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 64 53 25 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 59 55 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 64 53 59 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 55 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 51 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 64 45 51 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 35 27 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 48 46 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 64 53 48 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 34 26 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 24 25 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 43 36 64 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 64 24 43 64 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 23 62 22 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 22 61 63 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 23 59 61 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 23 60 21 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 21 56 58 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 23 55 20 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 20 53 57 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 23 62 19 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 19 52 54 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 23 51 52 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00049 23 62 18 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 18 49 50 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 23 48 49 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 23 46 17 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 17 45 47 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 23 44 60 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 23 43 16 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 16 63 44 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 23 55 15 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 15 45 42 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 23 41 56 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 23 46 14 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 14 53 40 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 23 54 13 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 13 50 41 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 23 36 12 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 12 37 38 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 23 35 11 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 11 34 39 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 23 40 33 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 23 36 10 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 10 31 32 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 23 62 36 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 23 62 9 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 9 30 29 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 23 42 30 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 23 62 8 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 8 33 28 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 23 47 31 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 23 38 7 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 7 32 27 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 23 29 6 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 6 28 26 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 23 57 37 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 23 53 45 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 23 46 5 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 5 53 25 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 23 55 4 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 4 53 59 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 23 46 55 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 23 46 3 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 3 45 51 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 23 27 35 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 23 46 2 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 2 53 48 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 23 26 34 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 23 25 24 23 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 23 36 1 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 1 24 43 23 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C42 23 23 8.91119e-13
C41 24 23 4.942e-14
C40 25 23 8.219e-14
C39 26 23 8.411e-14
C38 27 23 9.155e-14
C37 28 23 6.056e-14
C36 29 23 6.731e-14
C35 30 23 4.822e-14
C34 31 23 6.502e-14
C33 32 23 7.256e-14
C32 33 23 6.622e-14
C31 34 23 1.3366e-13
C30 35 23 1.2865e-13
C29 36 23 1.8859e-13
C28 37 23 9.622e-14
C27 38 23 1.1243e-13
C26 39 23 2.954e-14
C25 40 23 7.355e-14
C24 41 23 6.011e-14
C23 42 23 9.611e-14
C22 43 23 1.8227e-13
C21 44 23 5.411e-14
C20 45 23 2.4058e-13
C19 46 23 2.919e-13
C18 47 23 1.4915e-13
C17 48 23 1.9427e-13
C16 49 23 5.062e-14
C15 50 23 1.3088e-13
C14 51 23 1.9187e-13
C13 52 23 5.062e-14
C12 53 23 3.0519e-13
C11 54 23 1.1651e-13
C10 55 23 2.5651e-13
C9 56 23 1.2982e-13
C8 57 23 1.7171e-13
C7 58 23 2.954e-14
C6 59 23 2.1587e-13
C5 60 23 9.937e-14
C4 61 23 5.062e-14
C3 62 23 3.0462e-13
C2 63 23 1.2968e-13
C1 64 23 9.24999e-13
.ends somador_1bit_genlib_ocp_1_rows_roteado


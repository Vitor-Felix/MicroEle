* Spice description of na2_x1
* Spice driver version -1258236751
* Date ( dd/mm/yyyy hh:mm:ss ): 17/05/2012 at 17:28:57

* INTERF i0 i1 nq vdd vss 


.subckt na2_x1 2 3 5 1 6 
* NET 1 = vdd
* NET 2 = i0
* NET 3 = i1
* NET 5 = nq
* NET 6 = vss
Mtr_00004 1 3 5 1 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 5 2 1 1 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 4 3 5 6 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 6 2 4 6 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C6 1 6 1.168e-14
C5 2 6 2.405e-14
C4 3 6 2.33e-14
C2 5 6 2.086e-14
C1 6 6 1.168e-14
.ends na2_x1


*
* Curvas do diodo entre dreno e source com graal
*

* Circuit description

.include inversor_6.spi
.include inversor_6_gordo.spi
.include inversor_res_paralelos.spi

*V2 10 30 0V
*               
V2 10 30 pulse (0V 1.8V 1ns 1ps 1ps 1ns 2ns)
*  a vdd vss y 
X1 10 20 30  40 inversor_6
X2 40 20 30  41 inversor_6
X3 40 20 30  42 inversor_6
X4 40 20 30  43 inversor_6
X5 40 20 30  44 inversor_6
X6 10 20 30  45 inversor_6
X7 10 20 30  46 inversor_6_gordo
X8 46 20 30  47 inversor_6
X9 47 20 30  48 inversor_6
X10 48 20 30  49 inversor_6
X11 49 20 30  50 inversor_6
X12 10 20 30  51 inversor_6_gordo
X13 10 20 30  52 inversor_res_paralelos

v1 20 30 1.8V
v3 30 0 0V

* Auxiliar voltage source
* VAUX 10 20 DC 0

.model tp pmos level = 54
.model tn nmos level = 54
* Analysis

*.dc v2 0 1.8 0.001
.tran 0.0001 3ns
.end

*
* Curvas do diodo entre dreno e source com graal
*

* Circuit description

.include inversor_novo.spi

V2 10 30 0V


*  a vdd vss y 
X1 10 20 30  40 inversor_novo

v1 20 30 1.8V
v3 30 0 0V

.model tp pmos level = 54
.model tn nmos level = 54
* Analysis

.dc v2 0 1.8 0.001
*.tran 0.0001 3ns
.end

* Spice description of somador_4bit_genlib_ocp_nero
* Spice driver version 270587057
* Date ( dd/mm/yyyy hh:mm:ss ): 13/08/2013 at  9:13:12

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] c_0 c_4 s[0] s[1] s[2] s[3] 
* INTERF vdd vss 


.subckt somador_4bit_genlib_ocp_nero 127 136 160 154 132 87 163 149 129 56 73 
+ 79 15 114 167 124 
* NET 15 = s[2]
* NET 22 = somador_0.snand10
* NET 23 = somador_0.snand11
* NET 27 = somador_1.snand12
* NET 28 = somador_1.snand13
* NET 30 = somador_1.snand15
* NET 32 = somador_1.snand11
* NET 34 = somador_1.snand17
* NET 36 = somador_1.snand14
* NET 37 = somador_1.snand16
* NET 40 = somador_2.snand12
* NET 41 = somador_2.snand13
* NET 45 = somador_2.snand1
* NET 47 = somador_0.snand1
* NET 48 = somador_0.snand2
* NET 49 = somador_0.snand14
* NET 50 = somador_0.snand16
* NET 51 = somador_1.sinv1
* NET 52 = somador_1.snand1
* NET 53 = somador_1.snand5
* NET 54 = somador_1.snand2
* NET 55 = somador_3.snand16
* NET 56 = c_4
* NET 57 = somador_2.snand5
* NET 58 = somador_2.snand7
* NET 59 = somador_2.sinv1
* NET 60 = somador_2.snand15
* NET 61 = somador_2.snand3
* NET 62 = somador_2.snand2
* NET 63 = somador_0.snand5
* NET 66 = somador_0.sinv1
* NET 69 = somador_0.snand7
* NET 70 = somador_0.sinv2
* NET 71 = somador_0.sinv3
* NET 73 = s[0]
* NET 77 = somador_1.snand7
* NET 79 = s[1]
* NET 82 = somador_0.snand8
* NET 86 = c_1
* NET 87 = b[1]
* NET 88 = somador_1.snand10
* NET 93 = somador_3.snand10
* NET 95 = somador_3.snand14
* NET 102 = somador_3.snand17
* NET 104 = somador_3.snand5
* NET 108 = somador_2.snand6
* NET 110 = somador_2.snand8
* NET 112 = somador_3.snand7
* NET 114 = s[3]
* NET 118 = somador_2.snand4
* NET 120 = c_2
* NET 123 = somador_2.sinv2
* NET 124 = vss
* NET 126 = somador_0.snand12
* NET 127 = a[0]
* NET 128 = somador_0.snand13
* NET 129 = c_0
* NET 130 = somador_0.snand15
* NET 131 = somador_0.snand17
* NET 132 = b[0]
* NET 133 = somador_0.snand3
* NET 134 = somador_0.snand4
* NET 135 = somador_0.snand6
* NET 136 = a[1]
* NET 137 = somador_1.snand3
* NET 138 = somador_1.snand6
* NET 139 = somador_1.snand8
* NET 140 = somador_1.sinv3
* NET 141 = somador_1.sinv2
* NET 142 = somador_1.snand4
* NET 143 = somador_3.snand1
* NET 144 = somador_3.sinv2
* NET 145 = somador_3.snand2
* NET 146 = somador_3.sinv3
* NET 147 = somador_3.snand4
* NET 148 = somador_3.snand11
* NET 149 = b[3]
* NET 150 = somador_3.snand3
* NET 151 = somador_3.snand6
* NET 152 = somador_3.snand8
* NET 153 = somador_3.snand15
* NET 154 = a[3]
* NET 155 = somador_3.snand13
* NET 156 = somador_2.snand17
* NET 157 = somador_3.sinv1
* NET 158 = somador_3.snand12
* NET 159 = c_3
* NET 160 = a[2]
* NET 161 = somador_2.snand16
* NET 162 = somador_2.sinv3
* NET 163 = b[2]
* NET 164 = somador_2.snand11
* NET 165 = somador_2.snand10
* NET 166 = somador_2.snand14
* NET 167 = vdd
Mtr_00312 166 165 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 167 164 166 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 164 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 167 162 164 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 161 160 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 167 166 161 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 159 161 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00305 167 156 159 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 158 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 167 159 158 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 155 154 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 167 159 155 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 153 158 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 167 155 153 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 152 154 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 167 151 152 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 150 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 167 159 150 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 151 150 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 167 147 151 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 148 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 167 146 148 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 145 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 167 146 145 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 147 144 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 167 146 147 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 143 144 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 167 159 143 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 146 159 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 142 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 167 140 142 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 138 137 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 167 142 138 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 139 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 167 138 139 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 135 133 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 167 134 135 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 133 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 167 129 133 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 131 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 167 130 131 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 128 127 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 167 129 128 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 130 126 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 167 128 130 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 123 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 165 123 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 167 120 165 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 118 123 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 167 162 118 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 162 120 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 114 112 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 167 152 114 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 110 160 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 167 108 110 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 112 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 167 104 112 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 102 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 167 153 102 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 104 143 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 167 145 104 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 144 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 95 93 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 167 148 95 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 93 144 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 167 159 93 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 88 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 167 86 88 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 141 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 137 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 167 86 137 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 82 127 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00240 167 135 82 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00239 79 77 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 167 139 79 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 73 69 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 167 82 73 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 134 70 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 167 71 134 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 126 66 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 167 129 126 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 69 66 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 167 63 69 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 62 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 167 162 62 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 61 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 167 120 61 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 156 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 167 60 156 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 108 61 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 167 118 108 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 59 160 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 58 59 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 167 57 58 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 157 154 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 56 55 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 167 102 56 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 55 154 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 167 95 55 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 54 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 167 140 54 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 53 52 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 167 54 53 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 52 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 167 86 52 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 140 86 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 77 51 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 167 53 77 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 86 50 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 167 131 86 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 50 127 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 167 49 50 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 71 129 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 48 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 167 71 48 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 63 47 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 167 48 63 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 66 127 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 57 45 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 167 62 57 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 45 123 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 167 120 45 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 41 160 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 167 120 41 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 60 40 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 167 41 60 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 15 58 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 167 110 15 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 40 59 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 167 120 40 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 37 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 167 36 37 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 120 37 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 167 34 120 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 32 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 167 140 32 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 36 88 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 167 32 36 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 34 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 167 30 34 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 30 27 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 167 28 30 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 27 51 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 167 86 27 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 28 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 167 86 28 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 51 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 49 22 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 167 23 49 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 23 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 167 71 23 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 22 70 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 167 129 22 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 47 70 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 167 129 47 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 70 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 124 165 125 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 125 164 166 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 124 163 122 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 122 162 164 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 124 160 119 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 119 166 161 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 124 161 116 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 116 156 159 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 124 157 115 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 115 159 158 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 124 154 111 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 111 159 155 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 124 158 106 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 106 155 153 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 124 154 107 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 107 151 152 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 124 149 103 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 103 159 150 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 124 150 100 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 100 147 151 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 124 149 99 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 99 146 148 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 124 149 97 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 97 146 145 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 124 144 96 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 96 146 147 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 124 144 92 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 92 159 143 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 124 159 146 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 124 141 89 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 89 140 142 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 124 137 85 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 85 142 138 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 124 136 83 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 83 138 139 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 124 133 80 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 80 134 135 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 124 132 75 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 75 129 133 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 124 132 76 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 76 130 131 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 124 127 68 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 68 129 128 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 124 126 65 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 65 128 130 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 124 163 123 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00110 124 123 121 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 121 120 165 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 124 123 117 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 117 162 118 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 124 120 162 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 124 112 113 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 113 152 114 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 124 160 109 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 109 108 110 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 124 157 105 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 105 104 112 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 124 149 101 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 101 153 102 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 124 143 98 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 98 145 104 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 124 149 144 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00094 124 93 94 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 94 148 95 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 124 144 91 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 91 159 93 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 124 141 90 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 90 86 88 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 124 87 141 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 124 87 84 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 84 86 137 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 124 127 81 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 81 135 82 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 124 77 78 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 78 139 79 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 124 69 74 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 74 82 73 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 124 70 72 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 72 71 134 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 124 66 67 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 67 129 126 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 124 66 64 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 64 63 69 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 124 163 46 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 46 162 62 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 124 163 44 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 44 120 61 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 124 163 43 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 43 60 156 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 124 61 42 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 42 118 108 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 124 160 59 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 124 59 39 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 39 57 58 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 124 154 157 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00061 124 55 38 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 38 102 56 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 124 154 35 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 35 95 55 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 124 87 33 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 33 140 54 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 124 52 31 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 31 54 53 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 124 141 29 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 29 86 52 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 124 86 140 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00050 124 51 26 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 26 53 77 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 124 50 25 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 25 131 86 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 124 127 24 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 24 49 50 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 124 129 71 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 124 132 21 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 21 71 48 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 124 47 20 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 20 48 63 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 124 127 66 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 124 45 19 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 19 62 57 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 124 123 18 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 18 120 45 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 124 160 17 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 17 120 41 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 124 40 16 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 16 41 60 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 124 58 14 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 14 110 15 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 124 59 13 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 13 120 40 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 124 136 12 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 12 36 37 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 124 37 11 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 11 34 120 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 124 87 10 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 10 140 32 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 124 88 9 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 9 32 36 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 124 87 8 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 8 30 34 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 124 27 7 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 7 28 30 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 124 51 6 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 6 86 27 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 124 136 5 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 5 86 28 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 124 136 51 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 124 22 4 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 4 23 49 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 124 132 3 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 3 71 23 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 124 70 2 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 2 129 22 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 124 70 1 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 1 129 47 124 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 124 132 70 124 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C156 15 124 2.954e-14
C148 22 124 5.771e-14
C147 23 124 4.976e-14
C143 27 124 5.291e-14
C142 28 124 5.456e-14
C140 30 124 4.976e-14
C138 32 124 5.456e-14
C136 34 124 6.536e-14
C134 36 124 6.656e-14
C133 37 124 5.291e-14
C130 40 124 6.251e-14
C129 41 124 5.456e-14
C125 45 124 5.531e-14
C122 47 124 5.531e-14
C121 48 124 5.216e-14
C120 49 124 5.816e-14
C119 50 124 5.291e-14
C118 51 124 9.826e-14
C117 52 124 5.531e-14
C116 53 124 6.296e-14
C115 54 124 5.456e-14
C114 55 124 5.531e-14
C113 56 124 2.954e-14
C112 57 124 9.464e-14
C111 58 124 6.419e-14
C110 59 124 8.458e-14
C109 60 124 6.296e-14
C108 61 124 6.011e-14
C107 62 124 5.576e-14
C105 63 124 5.936e-14
C102 66 124 9.106e-14
C99 69 124 6.251e-14
C98 70 124 1.2787e-13
C97 71 124 1.2234e-13
C95 73 124 2.954e-14
C91 77 124 6.011e-14
C89 79 124 2.954e-14
C86 82 124 5.696e-14
C82 86 124 2.1737e-13
C81 87 124 1.8045e-13
C80 88 124 7.739e-14
C75 93 124 5.291e-14
C73 95 124 6.224e-14
C66 102 124 5.576e-14
C64 104 124 5.936e-14
C60 108 124 6.824e-14
C58 110 124 7.304e-14
C56 112 124 6.251e-14
C54 114 124 2.954e-14
C50 118 124 6.344e-14
C48 120 124 2.5609e-13
C45 123 124 1.4187e-13
C44 124 124 2.16836e-12
C42 126 124 5.771e-14
C41 127 124 1.6188e-13
C40 128 124 5.216e-14
C39 129 124 2.2343e-13
C38 130 124 5.456e-14
C37 131 124 7.784e-14
C36 132 124 1.9773e-13
C35 133 124 5.291e-14
C34 134 124 6.296e-14
C33 135 124 5.936e-14
C32 136 124 1.8372e-13
C31 137 124 5.531e-14
C30 138 124 5.216e-14
C29 139 124 6.416e-14
C28 140 124 1.5514e-13
C27 141 124 1.2427e-13
C26 142 124 5.216e-14
C25 143 124 7.427e-14
C24 144 124 1.1587e-13
C23 145 124 5.816e-14
C22 146 124 1.1074e-13
C21 147 124 5.936e-14
C20 148 124 6.656e-14
C19 149 124 1.6301e-13
C18 150 124 5.051e-14
C17 151 124 5.456e-14
C16 152 124 6.776e-14
C15 153 124 6.896e-14
C14 154 124 1.482e-13
C13 155 124 5.216e-14
C12 156 124 7.616e-14
C11 157 124 1.0906e-13
C10 158 124 5.531e-14
C9 159 124 2.3897e-13
C8 160 124 1.6764e-13
C7 161 124 5.291e-14
C6 162 124 1.4746e-13
C5 163 124 1.6917e-13
C4 164 124 5.216e-14
C3 165 124 6.131e-14
C2 166 124 6.176e-14
C1 167 124 2.23585e-12
.ends somador_4bit_genlib_ocp_nero


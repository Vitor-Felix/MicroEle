* Spice description of somador_4bit_genlib_4_rows_roteado
* Spice driver version 270587057
* Date ( dd/mm/yyyy hh:mm:ss ):  2/12/2014 at 15:19:22

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] c_0 c_4 s[0] s[1] s[2] s[3] 
* INTERF vdd vss 


.subckt somador_4bit_genlib_4_rows_roteado 204 177 225 220 197 171 239 209 194 
+ 215 200 2 241 230 247 165 
* NET 2 = s[1]
* NET 21 = somador_1.sinv4
* NET 24 = somador_1.snand15
* NET 26 = somador_0.snand14
* NET 29 = somador_0.snand2
* NET 31 = somador_0.sinv12
* NET 37 = somador_2.sinv14
* NET 38 = somador_2.sinv15
* NET 39 = somador_3.snand13
* NET 43 = somador_2.snand20
* NET 45 = somador_2.snand16
* NET 48 = somador_2.sinv10
* NET 50 = somador_2.snand2
* NET 52 = somador_1.snand7
* NET 53 = somador_1.snand8
* NET 54 = somador_1.snand13
* NET 55 = somador_1.snand5
* NET 56 = somador_1.sinv11
* NET 57 = somador_1.snand17
* NET 58 = somador_1.snand12
* NET 59 = somador_1.snand16
* NET 60 = somador_1.sinv10
* NET 61 = somador_0.sinv5
* NET 62 = somador_1.snand20
* NET 63 = somador_0.snand18
* NET 64 = somador_0.sinv3
* NET 65 = somador_0.snand3
* NET 66 = somador_0.sinv7
* NET 67 = somador_3.snand15
* NET 68 = somador_3.snand18
* NET 69 = somador_3.snand21
* NET 70 = somador_3.snand8
* NET 71 = somador_3.snand7
* NET 72 = somador_2.snand21
* NET 73 = somador_2.snand3
* NET 74 = somador_2.sinv2
* NET 75 = somador_2.sinv6
* NET 76 = somador_2.snand7
* NET 77 = somador_1.snand10
* NET 78 = somador_1.sinv9
* NET 80 = somador_1.sinv7
* NET 81 = somador_1.sinv13
* NET 82 = somador_1.snand14
* NET 86 = somador_1.sinv1
* NET 87 = somador_1.snand6
* NET 91 = somador_1.snand2
* NET 92 = somador_1.sinv5
* NET 98 = somador_0.sinv11
* NET 100 = somador_0.snand19
* NET 102 = somador_0.snand17
* NET 104 = somador_0.snand16
* NET 105 = somador_0.sinv10
* NET 109 = somador_0.snand13
* NET 112 = somador_0.snand12
* NET 115 = somador_0.sinv2
* NET 118 = somador_3.sinv13
* NET 119 = somador_3.snand19
* NET 122 = somador_3.snand14
* NET 123 = somador_3.sinv12
* NET 126 = somador_3.sinv3
* NET 131 = somador_3.snand16
* NET 134 = somador_3.snand20
* NET 135 = somador_3.snand3
* NET 136 = somador_3.sinv6
* NET 138 = somador_3.sinv2
* NET 139 = somador_3.sinv7
* NET 142 = somador_3.snand1
* NET 144 = somador_2.snand19
* NET 146 = somador_3.snand10
* NET 147 = somador_2.snand12
* NET 150 = somador_2.snand17
* NET 151 = somador_2.sinv13
* NET 154 = somador_2.snand4
* NET 156 = somador_2.sinv5
* NET 161 = somador_2.sinv7
* NET 163 = somador_2.snand8
* NET 164 = somador_2.snand10
* NET 165 = vss
* NET 167 = somador_1.sinv3
* NET 168 = somador_1.snand3
* NET 169 = somador_1.sinv6
* NET 170 = somador_1.sinv2
* NET 171 = b[1]
* NET 172 = c_1
* NET 173 = somador_1.snand4
* NET 174 = somador_1.snand1
* NET 175 = somador_1.sinv12
* NET 176 = somador_1.snand9
* NET 177 = a[1]
* NET 178 = somador_1.sinv8
* NET 179 = somador_1.snand19
* NET 180 = somador_1.snand21
* NET 181 = somador_0.snand20
* NET 182 = somador_1.snand18
* NET 183 = somador_1.sinv15
* NET 184 = somador_0.sinv14
* NET 185 = somador_0.snand15
* NET 186 = somador_1.sinv14
* NET 187 = somador_0.sinv13
* NET 188 = somador_0.snand21
* NET 189 = somador_0.snand6
* NET 190 = somador_0.sinv15
* NET 191 = somador_0.snand9
* NET 192 = somador_0.sinv1
* NET 193 = somador_0.snand5
* NET 194 = c_0
* NET 195 = somador_0.sinv9
* NET 196 = somador_0.snand4
* NET 197 = b[0]
* NET 198 = somador_0.sinv8
* NET 199 = somador_0.snand1
* NET 200 = s[0]
* NET 201 = somador_0.sinv4
* NET 202 = somador_0.snand8
* NET 203 = somador_0.snand10
* NET 204 = a[0]
* NET 205 = somador_0.snand7
* NET 206 = somador_3.sinv10
* NET 207 = somador_0.sinv6
* NET 208 = somador_3.snand12
* NET 209 = b[3]
* NET 210 = c_3
* NET 211 = somador_3.snand4
* NET 212 = somador_3.snand2
* NET 213 = somador_3.sinv5
* NET 214 = somador_3.sinv14
* NET 215 = c_4
* NET 216 = somador_3.snand17
* NET 217 = somador_3.sinv11
* NET 218 = somador_3.sinv15
* NET 219 = somador_3.sinv4
* NET 220 = a[3]
* NET 221 = somador_3.snand6
* NET 222 = somador_3.snand5
* NET 223 = somador_3.sinv1
* NET 224 = somador_3.snand9
* NET 225 = a[2]
* NET 226 = somador_2.snand18
* NET 227 = somador_3.sinv9
* NET 228 = c_2
* NET 229 = somador_3.sinv8
* NET 230 = s[3]
* NET 231 = somador_2.snand13
* NET 232 = somador_2.snand15
* NET 233 = somador_2.sinv12
* NET 234 = somador_2.sinv11
* NET 235 = somador_2.snand1
* NET 236 = somador_2.sinv4
* NET 237 = somador_2.sinv1
* NET 238 = somador_2.sinv3
* NET 239 = b[2]
* NET 240 = somador_2.snand14
* NET 241 = s[2]
* NET 242 = somador_2.sinv8
* NET 243 = somador_2.sinv9
* NET 244 = somador_2.snand6
* NET 245 = somador_2.snand5
* NET 246 = somador_2.snand9
* NET 247 = vdd
Mtr_00472 246 245 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 247 244 246 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 242 246 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00469 241 242 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00468 247 243 241 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00467 240 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 247 238 240 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00465 245 237 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 247 236 245 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 236 235 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00462 233 240 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 234 231 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 232 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00459 247 228 232 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00458 230 229 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00457 247 227 230 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00456 229 224 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00455 226 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00454 247 233 226 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00453 224 222 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 247 221 224 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 223 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00450 222 223 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00449 247 219 222 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 216 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 247 217 216 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00446 215 214 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00445 247 218 215 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00444 221 223 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00443 247 213 221 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 213 212 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 211 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 247 210 211 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 206 208 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00438 205 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00437 247 207 205 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00436 203 205 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00435 247 202 203 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 208 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00433 247 210 208 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00432 201 199 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00431 200 198 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00430 247 195 200 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00429 196 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00428 247 194 196 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00427 198 191 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 193 192 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 247 201 193 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00424 191 193 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 247 189 191 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 190 188 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 187 185 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 228 186 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 247 183 228 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00418 184 181 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00417 180 182 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00416 247 179 180 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00415 183 180 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00414 178 176 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00413 182 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00412 247 175 182 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00411 173 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00410 247 172 173 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00409 174 170 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00408 247 172 174 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 169 168 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 168 170 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 247 167 168 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 243 164 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 163 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 247 161 163 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00401 244 237 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 247 156 244 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00399 154 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 247 228 154 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00397 161 154 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00396 237 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00395 150 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00394 247 234 150 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00393 151 232 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00392 147 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00391 247 228 147 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 227 146 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 144 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00388 247 151 144 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00387 219 142 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00386 139 211 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 142 138 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 247 210 142 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 136 135 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 214 134 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 131 223 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 247 206 131 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 134 131 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 247 216 134 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 135 138 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 247 126 135 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00375 123 122 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00374 119 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00373 247 118 119 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00372 122 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00371 247 126 122 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00370 115 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00369 195 203 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00368 199 115 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00367 247 194 199 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00366 112 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00365 247 194 112 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00364 109 115 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 247 194 109 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 104 192 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 247 105 104 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 105 112 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 102 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00358 247 98 102 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 100 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00356 247 187 100 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00355 181 104 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00354 247 102 181 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 172 184 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 247 190 172 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 167 172 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 91 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00349 247 167 91 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00348 92 91 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00347 87 86 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 247 92 87 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 179 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 247 81 179 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 82 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00342 247 167 82 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00341 175 82 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00340 80 173 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00339 78 77 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00338 164 76 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 247 163 164 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 76 225 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 247 75 76 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 235 74 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 247 228 235 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00332 73 74 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 247 238 73 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00330 231 74 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00329 247 228 231 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 74 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 238 228 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00326 72 226 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00325 247 144 72 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00324 71 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00323 247 136 71 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00322 146 71 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00321 247 70 146 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00320 218 69 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00319 69 68 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 247 119 69 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 68 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 247 123 68 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 118 67 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00314 202 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00313 247 66 202 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00312 212 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 247 126 212 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 65 115 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 247 64 65 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 66 196 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 98 109 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 192 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00305 188 63 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 247 100 188 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 189 192 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 247 61 189 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 186 62 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 60 58 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 59 86 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 247 60 59 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 62 59 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 247 57 62 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 57 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 247 56 57 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 176 55 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 247 87 176 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 56 54 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 54 170 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 247 172 54 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 53 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 247 80 53 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 52 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 247 169 52 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 156 50 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 75 73 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 45 237 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 247 48 45 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 50 239 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 247 238 50 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 43 45 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 247 150 43 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 48 147 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 37 43 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 38 72 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 70 220 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 247 139 70 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 210 37 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 247 38 210 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 217 39 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 39 138 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 247 210 39 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 138 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 67 209 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 247 210 67 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 207 65 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 126 210 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 185 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 247 194 185 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 64 194 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 29 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 247 64 29 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 26 197 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 247 64 26 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 63 204 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 247 31 63 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 61 29 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 58 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 247 172 58 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 31 26 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 24 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 247 172 24 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 81 24 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 86 177 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 55 86 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 247 21 55 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 170 171 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 21 174 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00240 77 52 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00239 247 53 77 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 2 178 247 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 247 78 2 247 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 165 245 166 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 166 244 246 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 165 246 242 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00233 165 242 160 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 160 243 241 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 165 239 158 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 158 238 240 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 165 237 155 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 155 236 245 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 165 235 236 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00226 165 240 233 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00225 165 231 234 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00224 165 239 152 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 152 228 232 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 165 229 148 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 148 227 230 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 165 224 229 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00219 165 225 145 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 145 233 226 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 165 222 141 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 141 221 224 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 165 220 223 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 165 223 137 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 137 219 222 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 165 220 133 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 133 217 216 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 165 214 132 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 132 218 215 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 165 223 129 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 129 213 221 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 165 212 213 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00205 165 209 125 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 125 210 211 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 165 208 206 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 165 204 121 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 121 207 205 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 165 205 117 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 117 202 203 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 165 209 116 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 116 210 208 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 165 199 201 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 165 198 113 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 113 195 200 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 165 197 110 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 110 194 196 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 165 191 198 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00190 165 192 106 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 106 201 193 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 165 193 103 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 103 189 191 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 165 188 190 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00185 165 185 187 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00184 165 186 97 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 97 183 228 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 165 181 184 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00181 165 182 94 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 94 179 180 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 165 180 183 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 165 176 178 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 165 177 89 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 89 175 182 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 165 171 85 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 85 172 173 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 165 170 84 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 84 172 174 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 165 168 169 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00170 165 170 79 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 79 167 168 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 165 164 243 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00167 165 225 162 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 162 161 163 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 165 237 159 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 159 156 244 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 165 239 157 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 157 228 154 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 165 154 161 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00160 165 225 237 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00159 165 225 153 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 153 234 150 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 165 232 151 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00156 165 239 149 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 149 228 147 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 165 146 227 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 165 225 143 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 143 151 144 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 165 142 219 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 165 211 139 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00149 165 138 140 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 140 210 142 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 165 135 136 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 165 134 214 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 165 223 130 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 130 206 131 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 165 131 128 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 128 216 134 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 165 138 127 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 127 126 135 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 165 122 123 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00138 165 220 124 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 124 118 119 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 165 209 120 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 120 126 122 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 165 197 115 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00133 165 203 195 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00132 165 115 114 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 114 194 199 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 165 197 111 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 111 194 112 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 165 115 108 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 108 194 109 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 165 192 107 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 107 105 104 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 165 112 105 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00123 165 204 101 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 101 98 102 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 165 204 99 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 99 187 100 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 165 104 96 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 96 102 181 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 165 184 95 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 95 190 172 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 165 172 167 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 165 171 93 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 93 167 91 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 165 91 92 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 165 86 90 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 90 92 87 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 165 177 88 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 88 81 179 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 165 171 83 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 83 167 82 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 165 82 175 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 165 173 80 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00103 165 77 78 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00102 165 76 51 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 51 163 164 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 165 225 49 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 49 75 76 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 165 74 47 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 47 228 235 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 165 74 46 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 46 238 73 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 165 74 44 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 44 228 231 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 165 239 74 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 165 228 238 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 165 226 42 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 42 144 72 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 165 220 41 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 41 136 71 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 165 71 40 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 40 70 146 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 165 69 218 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00083 165 68 36 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 36 119 69 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 165 220 35 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00080 35 123 68 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 165 67 118 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00078 165 204 34 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 34 66 202 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 165 209 33 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 33 126 212 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 165 115 32 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 32 64 65 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 165 196 66 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00071 165 109 98 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00070 165 204 192 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 165 63 30 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 30 100 188 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 165 192 28 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 28 61 189 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 165 62 186 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 165 58 60 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 165 86 27 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 27 60 59 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 165 59 25 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 25 57 62 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 165 177 23 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 23 56 57 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 165 55 22 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 22 87 176 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 165 54 56 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 165 170 20 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 20 172 54 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 165 177 19 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 19 80 53 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 165 177 18 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 18 169 52 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 165 50 156 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00047 165 73 75 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 165 237 17 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 17 48 45 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 165 239 16 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 16 238 50 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 165 45 15 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 15 150 43 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 165 147 48 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 165 43 37 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 165 72 38 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 165 220 14 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 14 139 70 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 165 37 13 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 13 38 210 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 165 39 217 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 165 138 12 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 12 210 39 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 165 209 138 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 165 209 11 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 11 210 67 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 165 65 207 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 165 210 126 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 165 197 10 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 10 194 185 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 165 194 64 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 165 197 9 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 9 64 29 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 165 197 8 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 8 64 26 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 165 204 7 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 7 31 63 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 165 29 61 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 165 171 6 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 6 172 58 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 165 26 31 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 165 171 5 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 5 172 24 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 165 24 81 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 165 177 86 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 165 86 4 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 4 21 55 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 165 171 170 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 165 174 21 165 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 165 52 3 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 3 53 77 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 165 178 1 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 1 78 2 165 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C249 2 165 2.954e-14
C229 21 165 5.182e-14
C226 24 165 5.051e-14
C224 26 165 7.331e-14
C221 29 165 6.731e-14
C219 31 165 6.382e-14
C213 37 165 6.337e-14
C212 38 165 5.902e-14
C211 39 165 5.411e-14
C207 43 165 5.891e-14
C205 45 165 6.011e-14
C202 48 165 6.502e-14
C200 50 165 6.731e-14
C197 52 165 6.011e-14
C196 53 165 5.576e-14
C195 54 165 5.171e-14
C194 55 165 5.651e-14
C193 56 165 5.302e-14
C192 57 165 4.976e-14
C191 58 165 5.891e-14
C190 59 165 5.051e-14
C189 60 165 4.942e-14
C188 61 165 5.782e-14
C187 62 165 6.011e-14
C186 63 165 5.651e-14
C185 64 165 1.1674e-13
C184 65 165 7.331e-14
C183 66 165 6.502e-14
C182 67 165 5.771e-14
C181 68 165 5.531e-14
C180 69 165 5.411e-14
C179 70 165 6.656e-14
C178 71 165 5.291e-14
C177 72 165 5.771e-14
C176 73 165 7.091e-14
C175 74 165 1.1779e-13
C174 75 165 5.542e-14
C173 76 165 5.531e-14
C171 77 165 7.787e-14
C170 78 165 6.454e-14
C168 80 165 5.302e-14
C167 81 165 7.39e-14
C166 82 165 5.051e-14
C162 86 165 1.3867e-13
C161 87 165 5.696e-14
C157 91 165 5.051e-14
C156 92 165 4.942e-14
C150 98 165 6.502e-14
C148 100 165 5.696e-14
C146 102 165 5.696e-14
C144 104 165 6.371e-14
C143 105 165 4.822e-14
C139 109 165 5.363e-14
C136 112 165 6.011e-14
C133 115 165 1.2499e-13
C130 118 165 5.902e-14
C129 119 165 7.832e-14
C126 122 165 5.651e-14
C125 123 165 6.19e-14
C122 126 165 1.3746e-13
C117 131 165 5.051e-14
C114 134 165 5.651e-14
C113 135 165 6.491e-14
C112 136 165 6.742e-14
C110 138 165 1.5019e-13
C109 139 165 7.75e-14
C106 142 165 5.531e-14
C104 144 165 5.816e-14
C102 146 165 7.139e-14
C101 147 165 8.339e-14
C98 150 165 7.616e-14
C97 151 165 5.782e-14
C94 154 165 5.291e-14
C92 156 165 7.942e-14
C87 161 165 6.502e-14
C85 163 165 5.936e-14
C84 164 165 5.651e-14
C83 165 165 3.57304e-12
C81 167 165 1.3762e-13
C80 168 165 5.171e-14
C79 169 165 7.03e-14
C78 170 165 1.4203e-13
C77 171 165 2.459e-13
C76 172 165 2.8305e-13
C75 173 165 6.371e-14
C74 174 165 8.171e-14
C73 175 165 6.382e-14
C72 176 165 7.331e-14
C71 177 165 2.3078e-13
C70 178 165 1.0153e-13
C69 179 165 6.824e-14
C68 180 165 5.051e-14
C67 181 165 6.179e-14
C66 182 165 6.011e-14
C65 183 165 5.662e-14
C64 184 165 5.737e-14
C63 185 165 1.2131e-13
C62 186 165 6.865e-14
C61 187 165 5.782e-14
C60 188 165 7.091e-14
C59 189 165 7.136e-14
C58 190 165 6.55e-14
C57 191 165 5.651e-14
C56 192 165 1.4179e-13
C55 193 165 5.051e-14
C54 194 165 2.0735e-13
C53 195 165 6.382e-14
C52 196 165 7.451e-14
C51 197 165 2.2694e-13
C50 198 165 5.617e-14
C49 199 165 5.531e-14
C48 200 165 2.954e-14
C47 201 165 6.262e-14
C46 202 165 7.904e-14
C45 203 165 5.651e-14
C44 204 165 2.5382e-13
C43 205 165 5.051e-14
C42 206 165 7.342e-14
C41 207 165 8.782e-14
C40 208 165 6.131e-14
C39 209 165 2.3046e-13
C38 210 165 2.8609e-13
C37 211 165 8.939e-14
C36 212 165 8.411e-14
C35 213 165 4.822e-14
C34 214 165 5.617e-14
C33 215 165 2.954e-14
C32 216 165 6.536e-14
C31 217 165 9.022e-14
C30 218 165 7.942e-14
C29 219 165 6.622e-14
C28 220 165 2.6726e-13
C27 221 165 6.776e-14
C26 222 165 5.651e-14
C25 223 165 1.2931e-13
C24 224 165 5.651e-14
C23 225 165 2.467e-13
C22 226 165 7.619e-14
C21 227 165 5.422e-14
C20 228 165 3.7817e-13
C19 229 165 5.137e-14
C18 230 165 2.954e-14
C17 231 165 7.691e-14
C16 232 165 5.651e-14
C15 233 165 6.622e-14
C14 234 165 5.422e-14
C13 235 165 8.459e-14
C12 236 165 4.822e-14
C11 237 165 1.6579e-13
C10 238 165 1.5642e-13
C9 239 165 2.4606e-13
C8 240 165 6.131e-14
C7 241 165 2.954e-14
C6 242 165 5.017e-14
C5 243 165 6.862e-14
C4 244 165 6.656e-14
C3 245 165 7.571e-14
C2 246 165 5.291e-14
C1 247 165 3.71248e-12
.ends somador_4bit_genlib_4_rows_roteado


* Spice description of inverso_cmos_2
* Spice driver version 270587057
* Date ( dd/mm/yyyy hh:mm:ss ): 26/10/2015 at 16:43:20

* INTERF a vdd vss y 


.subckt inverso_cmos_2 1 2 4 3 
* NET 1 = a
* NET 2 = vdd
* NET 3 = y
* NET 4 = vss
Mtr_00002 3 1 2 2 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 4 1 3 4 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
C4 1 4 1.667e-14
C3 2 4 9.03e-15
C2 3 4 1.003e-14
C1 4 4 9.03e-15
.ends inverso_cmos_2


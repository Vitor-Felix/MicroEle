
 
.include somador_4bit_genlib_4_rows_roteado.spi
.model tp pmos level=54
.model tn nmos level=54

* a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] c_0 c_4 s[0] s[1] s[2] s[3] vdd vss 


x1 10 11 12 13 20 21 22 23 30 40 50 51 52 53 60 70  somador_4bit_genlib_4_rows_roteado


v1 10 70 pulse(0 1.8V 40ns 1ps 1ps 40ns 80ns)
v2 11 70 pulse(0 1.8V 40ns 1ps 1ps 40ns 80ns)
v3 12 70 pulse(0 1.8V 40ns 1ps 1ps 40ns 80ns)
v4 13 70 pulse(0 1.8V 40ns 1ps 1ps 40ns 80ns)
v5 20 70 pulse(0 1.8V 80ns 1ps 1ps 80ns 160ns)
v6 21 70 pulse(0 1.8V 80ns 1ps 1ps 80ns 160ns)
v7 22 70 pulse(0 1.8V 80ns 1ps 1ps 80ns 160ns)
v8 23 70 pulse(0 1.8V 80ns 1ps 1ps 80ns 160ns)
v9 30 70 pulse(0 1.8V 20ns 1ps 1ps 20ns 40ns)

v11 60 70 1.8V
v12 70 0 0V
.tran 0.01 160ns
.end


* Spice description of inversor_1
* Spice driver version -63871863
* Date ( dd/mm/yyyy hh:mm:ss ): 16/10/2014 at 15:15:50

* INTERF vdd vss x y 


.subckt inversor_1 2 3 1 4 
* NET 1 = x
* NET 2 = vdd
* NET 3 = vss
* NET 4 = y
Mtr_00002 4 1 2 2 tp L=1U W=1U AS=2P AD=2P PS=6U PD=6U 
Mtr_00001 4 1 3 3 tn L=1U W=1U AS=2P AD=2P PS=6U PD=6U 
C4 1 3 1.727e-14
C3 2 3 9.03e-15
C2 3 3 9.03e-15
C1 4 3 1.003e-14
.ends inversor_1


*
* Curvas estáticas do inversor_1

* Circuit description

.include inversor_6.spi
.include inversor_6_gordo.spi


V1 20 30 1.8V
v2 10 30 0V DC

*   a vdd vss y 

 
X1 10 20 30 40 inversor_6
X2 10 20 30 41 inversor_6
X3 41 20 30 42 inversor_6
X4 42 20 30 43 inversor_6
X5 10 20 30 44 inversor_6_gordo

V3 30 0 DC 0

.model tp pmos level = 54
.model tn nmos level = 54

* Analysis

.dc v2 0.7 1.1 0.001
.end

* Spice description of somador_1bit_nero
* Spice driver version -1258236751
* Date ( dd/mm/yyyy hh:mm:ss ): 22/05/2012 at 17:45:19

* INTERF a b c cout s vdd vss 


.subckt somador_1bit_nero 27 39 41 33 9 44 24 
* NET 3 = snand13
* NET 7 = snand8
* NET 9 = s
* NET 13 = snand6
* NET 16 = snand3
* NET 19 = snand4
* NET 24 = vss
* NET 26 = snand12
* NET 27 = a
* NET 28 = snand15
* NET 29 = sinv1
* NET 30 = snand7
* NET 31 = snand17
* NET 32 = snand16
* NET 33 = cout
* NET 34 = snand11
* NET 35 = snand14
* NET 36 = snand10
* NET 37 = snand5
* NET 38 = sinv3
* NET 39 = b
* NET 40 = snand2
* NET 41 = c
* NET 42 = sinv2
* NET 43 = snand1
* NET 44 = vdd
Mtr_00078 43 42 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 44 41 43 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 40 39 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 44 38 40 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 37 43 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 44 40 37 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 36 42 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 44 41 36 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 35 36 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 44 34 35 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 33 32 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 44 31 33 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 31 39 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 44 28 31 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 30 29 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 44 37 30 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 32 27 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 44 35 32 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 29 27 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 26 29 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 44 41 26 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 42 39 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 38 41 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 34 39 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 44 38 34 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 19 42 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 44 38 19 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 16 39 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 44 41 16 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 13 16 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 44 19 13 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 9 30 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 44 7 9 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 7 27 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 44 13 7 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 28 26 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 44 3 28 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 3 27 44 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 44 41 3 44 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 24 42 25 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 25 41 43 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 24 39 23 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 23 38 40 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 24 43 21 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 21 40 37 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 24 42 18 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 18 41 36 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 24 36 17 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 17 34 35 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 24 32 14 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 14 31 33 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 24 39 10 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 10 28 31 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 24 29 11 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 11 37 30 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 24 27 6 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 6 35 32 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 24 27 29 24 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 24 29 2 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 2 41 26 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 24 39 42 24 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 24 41 38 24 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 24 39 22 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 22 38 34 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 24 42 20 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 20 38 19 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 24 39 15 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 15 41 16 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 24 16 12 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 12 19 13 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 24 30 8 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 8 7 9 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 24 27 5 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 5 13 7 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 24 26 4 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 4 3 28 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 24 27 1 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 1 41 3 24 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C42 3 24 4.976e-14
C38 7 24 4.976e-14
C36 9 24 2.954e-14
C32 13 24 5.816e-14
C29 16 24 5.291e-14
C26 19 24 6.176e-14
C21 24 24 5.5216e-13
C19 26 24 6.011e-14
C18 27 24 1.3068e-13
C17 28 24 6.776e-14
C16 29 24 8.338e-14
C15 30 24 5.651e-14
C14 31 24 4.976e-14
C13 32 24 6.251e-14
C12 33 24 2.954e-14
C11 34 24 7.016e-14
C10 35 24 6.656e-14
C9 36 24 5.051e-14
C8 37 24 7.376e-14
C7 38 24 1.225e-13
C6 39 24 1.9181e-13
C5 40 24 5.456e-14
C4 41 24 2.4943e-13
C3 42 24 1.4299e-13
C2 43 24 6.011e-14
C1 44 24 5.69521e-13
.ends somador_1bit_nero


* Spice description of somador_4bit_genlib_4rows_nero
* Spice driver version -1258236751
* Date ( dd/mm/yyyy hh:mm:ss ): 29/05/2012 at 17:35:15

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] c_0 c_4 s[0] s[1] s[2] s[3] 
* INTERF vdd vss 


.subckt somador_4bit_genlib_4rows_nero 72 87 153 163 134 146 94 157 129 
+ 18 73 78 110 166 167 127 
* NET 18 = c_4
* NET 21 = somador_0.snand11
* NET 23 = somador_0.snand14
* NET 27 = somador_0.snand16
* NET 28 = somador_0.snand17
* NET 30 = somador_1.snand15
* NET 33 = somador_1.snand12
* NET 34 = somador_1.snand13
* NET 38 = somador_2.snand17
* NET 40 = somador_2.snand14
* NET 41 = somador_2.snand16
* NET 45 = somador_3.snand16
* NET 48 = somador_0.snand3
* NET 49 = somador_0.snand13
* NET 50 = somador_0.snand15
* NET 51 = somador_0.snand12
* NET 52 = somador_1.snand6
* NET 53 = somador_1.snand3
* NET 54 = somador_2.snand2
* NET 55 = somador_2.snand1
* NET 56 = somador_2.snand10
* NET 57 = somador_3.snand14
* NET 58 = somador_3.snand10
* NET 59 = somador_3.snand11
* NET 60 = somador_3.snand13
* NET 61 = somador_3.snand15
* NET 62 = somador_3.snand17
* NET 64 = somador_0.snand6
* NET 66 = somador_0.snand10
* NET 71 = somador_0.snand8
* NET 72 = a[0]
* NET 73 = s[0]
* NET 76 = somador_1.snand8
* NET 78 = s[1]
* NET 81 = somador_1.snand7
* NET 83 = somador_1.sinv1
* NET 84 = somador_1.snand17
* NET 87 = a[1]
* NET 89 = somador_1.snand16
* NET 92 = somador_2.snand11
* NET 94 = b[2]
* NET 97 = somador_2.snand3
* NET 98 = somador_2.snand4
* NET 99 = somador_2.sinv2
* NET 100 = somador_2.sinv3
* NET 104 = somador_2.snand6
* NET 105 = somador_2.snand5
* NET 108 = somador_2.snand8
* NET 110 = s[2]
* NET 113 = somador_2.snand7
* NET 116 = somador_3.sinv3
* NET 118 = somador_3.snand2
* NET 122 = somador_3.snand5
* NET 124 = somador_3.snand12
* NET 127 = vss
* NET 128 = somador_0.snand4
* NET 129 = c_0
* NET 130 = somador_0.sinv2
* NET 131 = somador_0.sinv3
* NET 132 = somador_0.snand1
* NET 133 = somador_0.snand2
* NET 134 = b[0]
* NET 135 = somador_0.snand5
* NET 136 = somador_0.sinv1
* NET 137 = somador_0.snand7
* NET 138 = somador_1.snand2
* NET 139 = somador_1.snand1
* NET 140 = somador_1.snand5
* NET 141 = somador_1.sinv2
* NET 142 = somador_1.snand10
* NET 143 = somador_1.snand14
* NET 144 = somador_1.snand4
* NET 145 = c_1
* NET 146 = b[1]
* NET 147 = somador_1.snand11
* NET 148 = somador_1.sinv3
* NET 149 = somador_2.snand12
* NET 150 = somador_2.snand15
* NET 151 = somador_2.sinv1
* NET 152 = c_2
* NET 153 = a[2]
* NET 154 = somador_2.snand13
* NET 155 = somador_3.snand4
* NET 156 = somador_3.snand3
* NET 157 = b[3]
* NET 158 = c_3
* NET 159 = somador_3.sinv2
* NET 160 = somador_3.snand6
* NET 161 = somador_3.snand1
* NET 162 = somador_3.sinv1
* NET 163 = a[3]
* NET 164 = somador_3.snand8
* NET 165 = somador_3.snand7
* NET 166 = s[3]
* NET 167 = vdd
Mtr_00312 166 165 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 167 164 166 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 162 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 164 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00308 167 160 164 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 161 159 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 167 158 161 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00305 159 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 160 156 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 167 155 160 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00302 154 153 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 167 152 154 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00300 151 153 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00299 150 149 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00298 167 154 150 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00297 149 151 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00296 167 152 149 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 147 146 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 167 148 147 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 148 145 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 143 142 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 167 147 143 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 144 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 167 148 144 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 140 139 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 167 138 140 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00286 138 146 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 167 148 138 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 137 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00283 167 135 137 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00282 139 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00281 167 145 139 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 133 134 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00279 167 131 133 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 135 132 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 167 133 135 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 132 130 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 167 129 132 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 128 130 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 167 131 128 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00272 124 162 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00271 167 158 124 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00270 165 162 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00269 167 122 165 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 122 161 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 167 118 122 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00266 118 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00265 167 116 118 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00264 156 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00263 167 158 156 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 110 113 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 167 108 110 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 108 153 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 167 104 108 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 113 151 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 167 105 113 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 104 97 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 167 98 104 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 98 99 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 167 100 98 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 97 94 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00251 167 152 97 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00250 92 94 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00249 167 100 92 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00248 89 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00247 167 143 89 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00246 152 89 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00245 167 84 152 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 81 83 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 167 140 81 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00242 78 81 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00241 167 76 78 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00240 73 137 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00239 167 71 73 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 136 72 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 131 129 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 71 72 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 167 64 71 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 66 130 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 167 129 66 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00232 130 134 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 62 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 167 61 62 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 61 124 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 167 60 61 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 59 157 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 167 116 59 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 57 58 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 167 59 57 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 116 158 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00222 155 159 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00221 167 116 155 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 56 99 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 167 152 56 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 105 55 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 167 54 105 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 55 99 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00215 167 152 55 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 54 94 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 167 100 54 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 53 146 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 167 145 53 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 100 152 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00209 76 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00208 167 52 76 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 52 53 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 167 144 52 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 83 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 51 136 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 167 129 51 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 50 51 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 167 49 50 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 49 72 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 167 129 49 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 64 48 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 167 128 64 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00196 48 134 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00195 167 129 48 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 60 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 167 158 60 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 18 45 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 167 62 18 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 45 163 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00189 167 57 45 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 58 159 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 167 158 58 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00186 41 153 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 167 40 41 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 158 41 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 167 38 158 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 40 56 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 167 92 40 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00180 38 94 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00179 167 150 38 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 99 94 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 30 33 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 167 34 30 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 34 87 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 167 145 34 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00173 84 146 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00172 167 30 84 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 141 146 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 142 141 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 167 145 142 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 145 27 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 167 28 145 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 33 83 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 167 145 33 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 28 134 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 167 50 28 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 27 72 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 167 23 27 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 23 66 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 167 21 23 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 21 134 167 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 167 131 21 167 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 127 165 125 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 125 164 166 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 127 163 162 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 127 163 121 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 121 160 164 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00151 127 159 119 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00150 119 158 161 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 127 157 159 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 127 156 115 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 115 155 160 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 127 153 112 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 112 152 154 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 127 153 151 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 127 149 107 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 107 154 150 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 127 151 103 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 103 152 149 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00139 127 146 96 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 96 148 147 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 127 145 148 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00136 127 142 93 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00135 93 147 143 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00134 127 141 90 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 90 148 144 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 127 139 86 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 86 138 140 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 127 146 82 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 82 148 138 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 127 136 79 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 79 135 137 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 127 141 75 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 75 145 139 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 127 134 70 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 70 131 133 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 127 132 69 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00121 69 133 135 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 127 130 67 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 67 129 132 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 127 130 63 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 63 131 128 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 127 162 126 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 126 158 124 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 127 162 123 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 123 122 165 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 127 161 120 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 120 118 122 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 127 157 117 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 117 116 118 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 127 157 114 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 114 158 156 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 127 113 111 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00105 111 108 110 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00104 127 153 109 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 109 104 108 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 127 151 106 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 106 105 113 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 127 97 101 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00099 101 98 104 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00098 127 99 102 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00097 102 100 98 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 127 94 95 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 95 152 97 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 127 94 91 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00093 91 100 92 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00092 127 87 88 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 88 143 89 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 127 89 85 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 85 84 152 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 127 83 80 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 80 140 81 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00086 127 81 77 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00085 77 76 78 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00084 127 137 74 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 74 71 73 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 127 72 136 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 127 129 131 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 127 72 68 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 68 64 71 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 127 130 65 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 65 129 66 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 127 134 130 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 127 157 47 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 47 61 62 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 127 124 46 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 46 60 61 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 127 157 44 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 44 116 59 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 127 58 43 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 43 59 57 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 127 158 116 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00066 127 159 42 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 42 116 155 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 127 99 39 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00063 39 152 56 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00062 127 55 37 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 37 54 105 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00060 127 99 36 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00059 36 152 55 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 127 94 35 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 35 100 54 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 127 146 32 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 32 145 53 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 127 152 100 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00053 127 87 31 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 31 52 76 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 127 53 29 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 29 144 52 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 127 87 83 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00048 127 136 26 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 26 129 51 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00046 127 51 25 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 25 49 50 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 127 72 24 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 24 129 49 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 127 48 22 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 22 128 64 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 127 134 20 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 20 129 48 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 127 163 19 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 19 158 60 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 127 45 17 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 17 62 18 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 127 163 16 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 16 57 45 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 127 159 15 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 15 158 58 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 127 153 14 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 14 40 41 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00028 127 41 13 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 13 38 158 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 127 56 12 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 12 92 40 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 127 94 11 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 11 150 38 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 127 94 99 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 127 33 10 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 10 34 30 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 127 87 9 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 9 145 34 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 127 146 8 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 8 30 84 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 127 146 141 127 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 127 141 7 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 7 145 142 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 127 27 6 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 6 28 145 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 127 83 5 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 5 145 33 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 127 134 3 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 3 50 28 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 127 72 4 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 4 23 27 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00004 127 66 2 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 2 21 23 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 127 134 1 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 1 131 21 127 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C153 18 127 2.954e-14
C149 21 127 4.976e-14
C147 23 127 4.976e-14
C143 27 127 6.251e-14
C142 28 127 5.456e-14
C140 30 127 5.816e-14
C137 33 127 7.691e-14
C136 34 127 5.096e-14
C132 38 127 5.936e-14
C130 40 127 5.936e-14
C129 41 127 5.291e-14
C125 45 127 5.531e-14
C121 48 127 5.291e-14
C120 49 127 4.976e-14
C119 50 127 5.576e-14
C118 51 127 5.051e-14
C117 52 127 4.976e-14
C116 53 127 5.891e-14
C115 54 127 5.936e-14
C114 55 127 5.531e-14
C113 56 127 5.363e-14
C112 57 127 6.224e-14
C111 58 127 5.531e-14
C110 59 127 5.456e-14
C109 60 127 6.344e-14
C108 61 127 5.216e-14
C107 62 127 6.296e-14
C104 64 127 5.696e-14
C102 66 127 6.851e-14
C97 71 127 5.696e-14
C96 72 127 1.2828e-13
C95 73 127 2.954e-14
C92 76 127 6.176e-14
C90 78 127 2.954e-14
C87 81 127 5.051e-14
C85 83 127 1.0666e-13
C84 84 127 6.896e-14
C81 87 127 1.5132e-13
C79 89 127 5.051e-14
C76 92 127 9.464e-14
C74 94 127 1.6869e-13
C71 97 127 5.771e-14
C70 98 127 4.976e-14
C69 99 127 1.3411e-13
C68 100 127 1.2082e-13
C64 104 127 5.456e-14
C63 105 127 5.408e-14
C60 108 127 5.216e-14
C58 110 127 2.954e-14
C55 113 127 6.011e-14
C52 116 127 1.3602e-13
C50 118 127 5.216e-14
C46 122 127 5.216e-14
C44 124 127 6.131e-14
C41 127 127 2.16836e-12
C40 128 127 7.016e-14
C39 129 127 2.0615e-13
C38 130 127 1.1347e-13
C37 131 127 1.6402e-13
C36 132 127 5.291e-14
C35 133 127 5.216e-14
C34 134 127 2.0037e-13
C33 135 127 5.936e-14
C32 136 127 1.0162e-13
C31 137 127 5.651e-14
C30 138 127 4.976e-14
C29 139 127 6.251e-14
C28 140 127 5.936e-14
C27 141 127 1.6171e-13
C26 142 127 9.491e-14
C25 143 127 5.936e-14
C24 144 127 8.144e-14
C23 145 127 2.8377e-13
C22 146 127 1.9893e-13
C21 147 127 5.576e-14
C20 148 127 1.2234e-13
C19 149 127 5.291e-14
C18 150 127 7.976e-14
C17 151 127 9.178e-14
C16 152 127 2.7569e-13
C15 153 127 1.5708e-13
C14 154 127 5.696e-14
C13 155 127 6.608e-14
C12 156 127 5.771e-14
C11 157 127 1.7781e-13
C10 158 127 3.0033e-13
C9 159 127 1.5651e-13
C8 160 127 6.536e-14
C7 161 127 6.131e-14
C6 162 127 8.746e-14
C5 163 127 1.578e-13
C4 164 127 5.816e-14
C3 165 127 6.251e-14
C2 166 127 2.954e-14
C1 167 127 2.23584e-12
.ends somador_4bit_genlib_4rows_nero


*
* Curvas estáticas do inversor_1

* Circuit description

.include inversor_6.spi
.include inversor_6_gordo.spi

V1 20 30 1.8V
v2 10 30 0V DC

*   a vdd vss y  

X6 10 20 30 45 inversor_6
X7 10 20 30 46 inversor_6_gordo

V3 30 0 DC 0

.model tp pmos level = 54
.model tn nmos level = 54

* Analysis

.dc v2 0 1.8 0.001
.end

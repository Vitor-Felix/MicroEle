* Spice description of inv_x1
* Spice driver version -1258236751
* Date ( dd/mm/yyyy hh:mm:ss ): 17/05/2012 at 17:29:04

* INTERF i nq vdd vss 


.subckt inv_x1 1 3 2 4 
* NET 1 = i
* NET 2 = vdd
* NET 3 = nq
* NET 4 = vss
Mtr_00002 3 1 2 2 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 4 1 3 4 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C4 1 4 2.405e-14
C3 2 4 9.28e-15
C2 3 4 1.932e-14
C1 4 4 8.72e-15
.ends inv_x1

